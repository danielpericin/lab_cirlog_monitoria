CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 180 30 200 9
48 114 1872 1042
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 114 1872 1042
143654930 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 149 207 0 1 11
0 11
0
0 0 21104 0
2 0V
-6 -16 8 -8
3 SET
-43 -4 -22 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 149 342 0 1 11
0 12
0
0 0 21104 0
2 0V
-6 -16 8 -8
5 RESET
-58 -5 -23 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 150 279 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
5 CLOCK
-57 -5 -22 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
14 Logic Display~
6 892 296 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 874 296 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 855 296 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 838 296 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
5 4013~
219 475 297 0 6 22
0 11 4 13 12 4 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 FF3
-35 -63 -14 -55
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 2 0
1 U
3747 0 0
0
0
7 Ground~
168 496 530 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
7 74LS153
119 770 442 0 14 29
0 4 2 3 3 5 6 3 3 3
2 2 2 8 7
0
0 0 13040 0
7 74LS153
-24 -60 25 -52
4 MUX2
29 -66 57 -58
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
7 74LS153
119 563 442 0 14 29
0 3 2 4 4 5 6 4 4 4
2 2 2 10 9
0
0 0 13040 0
7 74LS153
-24 -60 25 -52
4 MUX1
30 -65 58 -57
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
5 4013~
219 357 297 0 6 22
0 11 13 15 12 13 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 FF2
-35 -64 -14 -56
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 2 1 0
1 U
8903 0 0
0
0
5 4013~
219 249 297 0 6 22
0 11 15 14 12 15 6
0
0 0 4720 0
4 4013
10 -60 38 -52
3 FF1
-32 -66 -11 -58
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 1 0
1 U
3834 0 0
0
0
41
0 0 3 0 0 4096 0 0 0 28 11 2
517 406
517 261
3 0 4 0 0 4096 0 11 0 0 29 2
531 424
505 424
6 6 6 0 0 12416 0 13 11 0 0 4
273 261
288 261
288 451
531 451
0 5 5 0 0 4224 0 0 10 5 0 4
405 361
729 361
729 442
738 442
6 5 5 0 0 0 0 12 11 0 0 4
381 261
405 261
405 442
531 442
10 0 2 0 0 4096 0 10 0 0 12 2
738 487
694 487
3 0 3 0 0 0 0 10 0 0 11 2
738 424
711 424
4 0 3 0 0 0 0 10 0 0 11 2
738 433
711 433
7 0 3 0 0 0 0 10 0 0 11 2
738 460
711 460
8 0 3 0 0 0 0 10 0 0 11 2
738 469
711 469
6 9 3 0 0 128 0 8 10 0 0 4
499 261
711 261
711 478
738 478
2 0 2 0 0 8192 0 10 0 0 19 3
738 415
694 415
694 512
5 1 4 0 0 4224 0 8 10 0 0 4
505 279
702 279
702 406
738 406
0 6 6 0 0 4240 0 0 10 3 0 4
288 370
720 370
720 451
738 451
1 14 7 0 0 4224 0 4 10 0 0 3
892 314
892 469
802 469
13 1 8 0 0 8320 0 10 5 0 0 3
802 424
874 424
874 314
14 1 9 0 0 12416 0 11 6 0 0 5
595 469
630 469
630 334
855 334
855 314
13 1 10 0 0 12416 0 11 7 0 0 5
595 424
622 424
622 324
838 324
838 314
12 0 2 0 0 8320 0 10 0 0 21 3
808 487
808 512
601 512
11 12 2 0 0 0 0 10 10 0 0 2
808 406
808 487
12 0 2 0 0 0 0 11 0 0 24 3
601 487
601 512
496 512
11 12 2 0 0 0 0 11 11 0 0 2
601 406
601 487
10 0 2 0 0 0 0 11 0 0 24 2
531 487
496 487
2 1 2 0 0 0 0 11 9 0 0 3
531 415
496 415
496 524
7 0 4 0 0 0 0 11 0 0 27 2
531 460
505 460
8 0 4 0 0 0 0 11 0 0 27 2
531 469
505 469
0 9 4 0 0 0 0 0 11 29 0 3
505 431
505 478
531 478
1 0 3 0 0 0 0 11 0 0 0 2
531 406
514 406
0 4 4 0 0 0 0 0 11 36 0 3
505 316
505 433
531 433
1 0 11 0 0 4096 0 13 0 0 32 2
249 240
249 207
1 0 11 0 0 0 0 12 0 0 32 2
357 240
357 207
1 1 11 0 0 4224 0 1 8 0 0 3
161 207
475 207
475 240
4 0 12 0 0 4096 0 13 0 0 35 2
249 303
249 342
4 0 12 0 0 0 0 12 0 0 35 2
357 303
357 342
1 4 12 0 0 4224 0 2 8 0 0 3
161 342
475 342
475 303
2 5 4 0 0 0 0 8 8 0 0 5
451 261
441 261
441 316
505 316
505 279
5 3 13 0 0 4224 0 12 8 0 0 2
387 279
451 279
1 3 14 0 0 4224 0 3 13 0 0 2
162 279
225 279
0 2 15 0 0 8320 0 0 13 41 0 5
280 279
280 314
216 314
216 261
225 261
5 2 13 0 0 0 0 12 12 0 0 5
387 279
387 316
324 316
324 261
333 261
5 3 15 0 0 0 0 13 12 0 0 2
279 279
333 279
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
